LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONDITIONCODEREGISTER IS
 PORT ( CLOCK, RESET,WRITEENABLE : IN STD_LOGIC;
 CCRIN : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
 CCROUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0) );
END CONDITIONCODEREGISTER; 

ARCHITECTURE BEHAVIOUR OF CONDITIONCODEREGISTER IS
 BEGIN
 PROCESS (CLOCK, RESET)
 BEGIN
IF RESET = '1' THEN 
CCROUT <= "0000";
ELSIF (RISING_EDGE(CLOCK)AND WRITEENABLE='1') THEN
CCROUT <= CCRIN;
END IF;
END PROCESS;
END BEHAVIOUR; 