LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DFF IS
PORT (D: IN STD_LOGIC;
	RST,CLK: IN STD_LOGIC;
	Q: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF DFF IS
BEGIN
	PROCESS (CLK,RST)
	BEGIN
		IF (RST='1') THEN
			Q <= '0';
		ELSIF (RISING_EDGE(CLK)) THEN
			Q <= D;
		END IF;
	END PROCESS;
END ARCHITECTURE;	


