LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DFF IS
Generic(N : integer := 32);
PORT (D: IN STD_LOGIC;
	RST,CLK: IN STD_LOGIC;
	Q: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF DFF IS
BEGIN
	PROCESS (CLK,RST)
	BEGIN
		IF (RISING_EDGE(CLK)) THEN
			IF (RST='1') THEN
				Q <= '0';
			ELSE 
				Q <= D;
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE;	

