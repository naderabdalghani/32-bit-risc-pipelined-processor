LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL; 
ENTITY DEC_EX_BUFFER IS PORT(
BUFFER_OUTPUT :OUT STD_LOGIC_VECTOR(131 DOWNTO 0);
READDATA1:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
READDATA:IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
EA: IN  STD_LOGIC_VECTOR(19 DOWNTO 0);
IMM:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
TWO_FETCHES:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
PREDICTION_SIGNAL:IN STD_LOGIC;
PC:IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
WRITE_REG1:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
WRITE_REG2:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
CLK:IN STD_LOGIC;
RST:IN STD_LOGIC;
BRANCH,MR,MW,P_IN,P_OUT,SP_INC,SP_DEC,CALL,WB1,WB2,RET,ALU_ENABLE,RTI,NO_OPERANDS,IGNORE_RSRC2: IN STD_LOGIC;
ALU_SELECTORS: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
OP_GROUP: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
READ_ADDRESS1_REGFILE,READ_ADDRESS2_REGFILE: IN STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END DEC_EX_BUFFER;
ARCHITECTURE BEHAVIORAL OF DEC_EX_BUFFER IS
SIGNAL READDATA2:STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

READDATA2 <= READDATA WHEN TWO_FETCHES ="00"
ELSE "000000000000" &EA WHEN TWO_FETCHES ="10"
ELSE STD_LOGIC_VECTOR(RESIZE(SIGNED(IMM), READDATA2'LENGTH))WHEN TWO_FETCHES ="01"
ELSE READDATA; 

 PROCESS(CLK,RST) 
 BEGIN
IF(RST='1'  ) THEN
BUFFER_OUTPUT <= (OTHERS => '0');

ELSIF(RISING_EDGE(CLK) ) THEN
BUFFER_OUTPUT <=  READ_ADDRESS1_REGFILE & READ_ADDRESS2_REGFILE & NO_OPERANDS & IGNORE_RSRC2 & BRANCH & MR & MW & P_IN & P_OUT & SP_INC &SP_DEC  & WB1 & WB2 & CALL & RET & ALU_ENABLE & RTI & ALU_SELECTORS & TWO_FETCHES & OP_GROUP & PREDICTION_SIGNAL & READDATA1 & READDATA2 & PC & WRITE_REG1 & WRITE_REG2;
END IF;


END PROCESS ;



END BEHAVIORAL ;
