LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DYNAMIC_BRANCH_ENABLE IS
PORT (BRANCHING_REG: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      WB1_CONTROL_UNIT, WB2_CONTROL_UNIT: IN STD_LOGIC;
      RDST_IF_ID ,RSRC_IF_ID: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      WB1_ID_EX ,WB2_ID_EX: IN STD_LOGIC;
      RDST_ID_EX ,RSRC_ID_EX: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      WB1_EX_MEM ,WB2_EX_MEM: IN STD_LOGIC;
      RDST_EX_MEM ,RSRC_EX_MEM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      WB1_MEM_WB ,WB2_MEM_WB: IN STD_LOGIC;
      RDST_MEM_WB ,RSRC_MEM_WB: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      ENABLE_DYNAMIC_PREDICTION: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE ARCH OF DYNAMIC_BRANCH_ENABLE IS
SIGNAL FIRST, SECOND, THIRD, FORTH: STD_LOGIC; -- SIGNAL IS '1' IF BRANCH WAITING FOR IT
SIGNAL FIRST1, FIRST2, SECOND1, SECOND2, THIRD1, THIRD2, FORTH1, FORTH2: STD_LOGIC;
SIGNAL SELECTOR11, SELECTOR12, SELECTOR21, SELECTOR22, SELECTOR31, SELECTOR32, SELECTOR41, SELECTOR42: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL REG11, REG12, REG21, REG22, REG31, REG32, REG41, REG42: STD_LOGIC_VECTOR(2 DOWNTO 0); -- SIGNAL IS '0' WHEN IT EQUALS TO BRANCHING REG
BEGIN
    -- IF ANY REG EQUALS TO "000" THEN IT'S THE SAME BRANCHING REGISTER
    REG11 <= RDST_IF_ID XOR BRANCHING_REG;
    REG12 <= RSRC_IF_ID XOR BRANCHING_REG;
    REG21 <= RDST_ID_EX XOR BRANCHING_REG;
    REG22 <= RSRC_ID_EX XOR BRANCHING_REG;
    REG31 <= RDST_EX_MEM XOR BRANCHING_REG;
    REG32 <= RSRC_EX_MEM XOR BRANCHING_REG;
    REG41 <= RDST_MEM_WB XOR BRANCHING_REG;
    REG42 <= RSRC_MEM_WB XOR BRANCHING_REG;

    -- SET SELECTORS
    SELECTOR11 <= REG11 & WB1_CONTROL_UNIT;
    SELECTOR12 <= REG12 & WB2_CONTROL_UNIT;
    SELECTOR21 <= REG21 & WB1_ID_EX;
    SELECTOR22 <= REG22 & WB2_ID_EX;
    SELECTOR31 <= REG31 & WB1_EX_MEM;
    SELECTOR32 <= REG32 & WB2_EX_MEM;
    SELECTOR41 <= REG41 & WB1_MEM_WB;
    SELECTOR42 <= REG42 & WB2_MEM_WB;

    WITH SELECTOR11 SELECT FIRST1 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;
    WITH SELECTOR12 SELECT FIRST2 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;

    WITH SELECTOR21 SELECT SECOND1 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;
    WITH SELECTOR22 SELECT SECOND2 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;

    WITH SELECTOR31 SELECT THIRD1 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;
    WITH SELECTOR32 SELECT THIRD2 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;

    WITH SELECTOR41 SELECT FORTH1 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;
    WITH SELECTOR42 SELECT FORTH2 <=
    '1' WHEN "0001",
    '0' WHEN OTHERS;


    -- SETTING SIGNALS TO CHECK IF BRANCH IS WAITING FOR ONE OF THEM
    FIRST <= FIRST1 OR FIRST2;
    SECOND <= SECOND1 OR SECOND2;
    THIRD <= THIRD1 OR THIRD2;
    FORTH <= FORTH1 OR FORTH2;


    ENABLE_DYNAMIC_PREDICTION <= NOT (FIRST OR SECOND OR THIRD OR FORTH);

END ARCHITECTURE;
