LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DFF IS
	GENERIC(N : INTEGER := 32);
	PORT (
		D: IN STD_LOGIC;
		RST,CLK: IN STD_LOGIC;
		Q: OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF DFF IS
BEGIN
	PROCESS (CLK,RST)
	BEGIN
		IF (RISING_EDGE(CLK)) THEN
			IF (RST='1') THEN
				Q <= '0';
			ELSE 
				Q <= D;
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE;
