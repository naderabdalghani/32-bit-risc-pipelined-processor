LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY REG IS
Generic(N : integer := 32);
PORT (D: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	RST,CLK,WR_ENABLE: IN STD_LOGIC;
	Q: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF REG IS
BEGIN
	PROCESS (CLK,RST)
	BEGIN
		IF (RISING_EDGE(CLK)) THEN
			IF (RST='1') THEN
				Q <= (OTHERS => '0');
			ELSIF (WR_ENABLE = '1') THEN
				Q <= D;
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE;	

