LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;

ENTITY DATA_MEMORY IS
	GENERIC (WORD_SIZE : INTEGER := 16; ADDRESS_WIDTH: INTEGER := 32; MEMORY_SIZE: INTEGER := 4096);
	PORT(	
		W  : IN STD_LOGIC;
		R  : IN STD_LOGIC;
		CLK  : IN STD_LOGIC;
		ADDRESS : IN  STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
		DATA_IN  : IN  STD_LOGIC_VECTOR(WORD_SIZE * 2 - 1 DOWNTO 0);
		DATA_OUT  : OUT  STD_LOGIC_VECTOR(WORD_SIZE * 2 - 1 DOWNTO 0));
END ENTITY DATA_MEMORY;

ARCHITECTURE BEHAVIORAL OF DATA_MEMORY IS
    TYPE MEMORY_TYPE IS ARRAY(MEMORY_SIZE - 1 DOWNTO 0) OF STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
    
	-- INPUT INSTRUCTION MEMORY DATA FROM ASSEMBLER PROGRAM OUTPUT

  	IMPURE FUNCTION FILL_MEMORY RETURN MEMORY_TYPE IS
		VARIABLE MEMORY_CONTENT : MEMORY_TYPE;
		VARIABLE TEXT_LINE : LINE;
		VARIABLE I: INTEGER;
        VARIABLE BINARY_TEXT_LINE : BIT_VECTOR(WORD_SIZE - 1 DOWNTO 0);
		FILE MEMORY_FILE: TEXT;
    BEGIN
        -- OPEN FILE
        FILE_OPEN(MEMORY_FILE, "MEM.OUT",  READ_MODE);

        -- STORE RESET PC ADDRESS & INTERRUPT PC ADDRESS
        I := 0;
        WHILE NOT ENDFILE(MEMORY_FILE) AND I < 4 LOOP
            READLINE(MEMORY_FILE, TEXT_LINE);
            READ(TEXT_LINE, BINARY_TEXT_LINE);
            -- REPORT "TEXT_LINE INSIDE MEMORY LOOP: "& INTEGER'IMAGE(TO_INTEGER(UNSIGNED(TO_STDLOGICVECTOR(BINARY_TEXT_LINE))));
            MEMORY_CONTENT(I) := TO_STDLOGICVECTOR(BINARY_TEXT_LINE);
            I := I + 1;
        END LOOP;

        FILE_CLOSE(MEMORY_FILE);
        RETURN MEMORY_CONTENT;

    END FUNCTION FILL_MEMORY;
    
    SIGNAL DATA_MEMORY : MEMORY_TYPE := FILL_MEMORY;

BEGIN
    PROCESS(CLK) IS
        BEGIN
        IF FALLING_EDGE(CLK) THEN
            IF W = '1' THEN
                DATA_MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))) <= DATA_IN(WORD_SIZE - 1 DOWNTO 0);
                DATA_MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 1) <= DATA_IN(WORD_SIZE * 2 - 1 DOWNTO WORD_SIZE);
            END IF;
            IF R = '1' THEN
                DATA_OUT <= DATA_MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 1) & DATA_MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)));    
            END IF ;
        END IF ;
    END PROCESS;
END BEHAVIORAL;