LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FETCHING_STAGE IS
PORT (DATA_EXE_STAGE, DATA_DATA_MEMORY: IN STD_LOGIC_VECTOR(31 DOWNTO 0);               
      WRONG_DECISION, LW_USE_CASE, INTERRUPT1, RETURN_INTERRUPT, RET: IN STD_LOGIC;     
      PC: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);                                            
      --------------------------- PC CIRCUIT I/O DONE --------------------------------
      INSTRUCTION_MEMORY: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      FE_ID: OUT STD_LOGIC_VECTOR(64 DOWNTO 0);
      TWO_FETCHES: OUT STD_LOGIC;
      -------------------------- FETCHING_CIRCUIT DONE -------------------------------
      WB1_CONTROL_UNIT, WB2_CONTROL_UNIT: IN STD_LOGIC;
      WB1_ID_EX ,WB2_ID_EX: IN STD_LOGIC;
      RDST_ID_EX ,RSRC_ID_EX: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      WB1_EX_MEM ,WB2_EX_MEM: IN STD_LOGIC;
      RDST_EX_MEM ,RSRC_EX_MEM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      WB1_MEM_WB ,WB2_MEM_WB: IN STD_LOGIC;
      RDST_MEM_WB ,RSRC_MEM_WB: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      ---------------------- ENABLE_DYNAMIC_PREDICTION DONE --------------------------
      DYNAMIC_BRANCH_ADDRESS: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      JUMPING_REG: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      JZ_EXE_STAGE,ZERO_FLAG: IN STD_LOGIC;
      BRANCHING_REG: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
      ---------------------- DYNAMIC_BRANCH_PREDICTION DONE --------------------------
      INTERRUPT_SIGNAL,RTI_SIGNAL_FROM_ALL_STAGES: IN STD_LOGIC;
      INT_TO_MEM_STAGE: OUT STD_LOGIC;
      ------------------------- INTERRUPT_HANDLER DONE -------------------------------
      CLK,RST: IN STD_LOGIC);
END ENTITY;

ARCHITECTURE ARCH OF FETCHING_STAGE IS
SIGNAL PC_SIGNAL: STD_LOGIC_VECTOR(31 DOWNTO 0); -- PC OUT
SIGNAL BRANCHING_REG_SIGNAL: STD_LOGIC_VECTOR(2 DOWNTO 0); -- TO GET THE REGISTER OF BRANCHING
SIGNAL TWO_FETCHES_BEFORE_DFF: STD_LOGIC; -- HOLDING TWO FETCHES SIGNAL BEFORE DFF
SIGNAL RDST_IF_ID ,RSRC_IF_ID: STD_LOGIC_VECTOR(2 DOWNTO 0); -- HOLDING RDST,RSRC FROM FE/ID BUFFER
SIGNAL FE_ID_SIGNAL: STD_LOGIC_VECTOR(64 DOWNTO 0); -- FE/ID SIGNAL
SIGNAL FIRST_16_BITS_INST_MEM: STD_LOGIC_VECTOR(15 DOWNTO 0); -- FIRST 16 BIT OF INSTRUCTION
SIGNAL ENABLE_DYNAMIC_PREDICTION: STD_LOGIC; -- ENABLE OF DYNAMIC BRANCH PREDICTION
SIGNAL PREDICTION_SIGNAL: STD_LOGIC; -- HOLDING PREDICTION SIGNAL FROM DYNAMIC BRANCH PREDICTION
SIGNAL PREDICTION_ADDRESS: STD_LOGIC_VECTOR(31 DOWNTO 0); -- ADDRESS TO BRANCH TO FROM DYNAMIC PREDICTION CIRCUIT
SIGNAL RESET_FETCHING_AND_STALL_PC: STD_LOGIC; -- TO STALL PC AND RESET FETCHING
BEGIN
    PC <= PC_SIGNAL;
    FE_ID <= FE_ID_SIGNAL;
    RDST_IF_ID <= FE_ID_SIGNAL(24 DOWNTO 22);
    RSRC_IF_ID <= FE_ID_SIGNAL(21 DOWNTO 19);
    BRANCHING_REG <= BRANCHING_REG_SIGNAL;
    TWO_FETCHES <= TWO_FETCHES_BEFORE_DFF;

    -- GETTING DATA FOR DYNAMIC BRANCH PREDICTION TEST
    WITH TWO_FETCHES_BEFORE_DFF SELECT BRANCHING_REG_SIGNAL <= -- GET RDST IN FIRST FETH ONLY (AS BRANCH IS A 16-BIT INSTRUCTION)
    INSTRUCTION_MEMORY(8 DOWNTO 6) WHEN '0',
    BRANCHING_REG_SIGNAL WHEN OTHERS;
    WITH TWO_FETCHES_BEFORE_DFF SELECT FIRST_16_BITS_INST_MEM <= -- GETTING THE FIRST 16-BIT OF THE INSTRUCTION
    INSTRUCTION_MEMORY WHEN '0',
    FIRST_16_BITS_INST_MEM WHEN OTHERS;


    -- PORT MAP PC CIRCUIT
    PC_CIRCUIT: ENTITY WORK.PC_CIRCUIT PORT MAP (DATA_EXE_STAGE, PREDICTION_ADDRESS, DATA_DATA_MEMORY ,CLK, RST, 
    WRONG_DECISION, PREDICTION_SIGNAL, RESET_FETCHING_AND_STALL_PC, LW_USE_CASE, INTERRUPT1, RETURN_INTERRUPT, RET,PC_SIGNAL);

    -- PORT MAP FETCHING BUFFER CIRCUIT
    FETCHING_CIRCUIT: ENTITY WORK.FETCHING_CIRCUIT PORT MAP (INSTRUCTION_MEMORY, PC_SIGNAL,
    RST, CLK, RESET_FETCHING_AND_STALL_PC, WRONG_DECISION, LW_USE_CASE, PREDICTION_SIGNAL, FE_ID_SIGNAL,TWO_FETCHES_BEFORE_DFF);

    -- PORT MAP DYNAMIC_PREDICTION_ENABLE
    DYNAMIC_PREDICTION_ENABLE: ENTITY WORK.DYNAMIC_BRANCH_ENABLE PORT MAP (BRANCHING_REG_SIGNAL,WB1_CONTROL_UNIT, WB2_CONTROL_UNIT,
    RDST_IF_ID ,RSRC_IF_ID,WB1_ID_EX ,WB2_ID_EX,RDST_ID_EX ,RSRC_ID_EX,WB1_EX_MEM ,WB2_EX_MEM,RDST_EX_MEM ,RSRC_EX_MEM,WB1_MEM_WB ,WB2_MEM_WB,
    RDST_MEM_WB ,RSRC_MEM_WB,ENABLE_DYNAMIC_PREDICTION);

    -- PORT MAP DYNAMIC BRANCH CIRCUIT
    DYNAMIC_BRANCH_PREDICTION: ENTITY WORK.DYNAMIC_BRANCH PORT MAP (DYNAMIC_BRANCH_ADDRESS, JUMPING_REG, FIRST_16_BITS_INST_MEM,
    ENABLE_DYNAMIC_PREDICTION, CLK, RST, JZ_EXE_STAGE, ZERO_FLAG, PREDICTION_SIGNAL, BRANCHING_REG_SIGNAL, PREDICTION_ADDRESS);

    -- PORT MAP INTERRUPT HANDLER
    INTERRUPT_HANDLER: ENTITY WORK.INT_HANDLER PORT MAP (INTERRUPT_SIGNAL, RTI_SIGNAL_FROM_ALL_STAGES, INTERRUPT1, CLK, RST, 
    INT_TO_MEM_STAGE, RESET_FETCHING_AND_STALL_PC);
END ARCHITECTURE;
