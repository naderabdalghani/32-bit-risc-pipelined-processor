LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY HAZARDDETECTION IS PORT (
LOAD:OUT STD_LOGIC;
DEC_EX_MEMREAD:IN STD_LOGIC;
F_DEC_SRC1,F_DEC_SRC2,DEC_EX_DEST:IN STD_LOGIC_VECTOR(2 DOWNTO 0) ;
OP_CODE:IN STD_LOGIC_VECTOR(6 DOWNTO 0);
NO_OPERANDS,IGNORE_RSRC2:IN STD_LOGIC;
TWO_FETCHES:IN STD_LOGIC
);
END HAZARDDETECTION ;
ARCHITECTURE BEHAVIORAL OF HAZARDDETECTION IS
    SIGNAL NO_OPERAND: STD_LOGIC;
BEGIN
    WITH OP_CODE SELECT NO_OPERAND <=
    '1' WHEN "0000000" | "0100111" | "0100101",
    '0' WHEN OTHERS;

LOAD <= '1' 
WHEN ( (
(F_DEC_SRC1 = DEC_EX_DEST  AND NO_OPERAND='0')
OR (F_DEC_SRC2 = DEC_EX_DEST  AND NO_OPERAND='0' AND IGNORE_RSRC2='0')
) 
AND DEC_EX_MEMREAD = '1' AND TWO_FETCHES = '0')
ELSE '0';



END BEHAVIORAL ;
