LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;

ENTITY INSTRUCTION_MEMORY IS
	GENERIC (WORD_SIZE : INTEGER := 16; ADDRESS_WIDTH: INTEGER := 32; MEMORY_SIZE: INTEGER := 4096);
	PORT(	
		CLK  : IN STD_LOGIC;
		WR  : IN STD_LOGIC;
		ADDRESS : IN  STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
		DATA_IN  : IN  STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
		DATA_OUT  : OUT  STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0));
END ENTITY INSTRUCTION_MEMORY;

ARCHITECTURE BEHAVIORAL OF INSTRUCTION_MEMORY IS
    TYPE MEMORY_TYPE IS ARRAY(MEMORY_SIZE - 1 DOWNTO 0) OF STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
    
	-- INPUT INSTRUCTION MEMORY DATA FROM ASSEMBLER PROGRAM OUTPUT

  	IMPURE FUNCTION FILL_MEMORY RETURN MEMORY_TYPE IS
		VARIABLE MEMORY_CONTENT : MEMORY_TYPE;
		VARIABLE TEXT_LINE : LINE;
		VARIABLE COUNT: INTEGER;
		VARIABLE I: INTEGER;
        VARIABLE STARTING_ADDRESS: STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
        VARIABLE BINARY_TEXT_LINE : BIT_VECTOR(WORD_SIZE - 1 DOWNTO 0);
		FILE MEMORY_FILE: TEXT;
    BEGIN
        -- OPEN FILE
        FILE_OPEN(MEMORY_FILE, "mem.out",  READ_MODE);

        -- READ FIRST 16 BITS OF STARTING ADDRESS
        READLINE(MEMORY_FILE, TEXT_LINE);
        READ(TEXT_LINE, BINARY_TEXT_LINE);
	    -- REPORT "TEXT_LINE: "& INTEGER'IMAGE(TO_INTEGER(UNSIGNED(TO_STDLOGICVECTOR(BINARY_TEXT_LINE))));
        STARTING_ADDRESS(WORD_SIZE - 1 DOWNTO 0) := TO_STDLOGICVECTOR(BINARY_TEXT_LINE); 

        -- READ SECOND 16 BITS OF STARTING ADDRESS
        READLINE(MEMORY_FILE, TEXT_LINE);
        READ(TEXT_LINE, BINARY_TEXT_LINE);
	    -- REPORT "TEXT_LINE: "& INTEGER'IMAGE(TO_INTEGER(UNSIGNED(TO_STDLOGICVECTOR(BINARY_TEXT_LINE))));
        STARTING_ADDRESS(ADDRESS_WIDTH - 1 DOWNTO WORD_SIZE) := TO_STDLOGICVECTOR(BINARY_TEXT_LINE); 

        COUNT := TO_INTEGER(UNSIGNED(STARTING_ADDRESS));

        -- SKIP INSTRUCTIONS UNTIL STARTING ADDRESS
        I := 0;
        WHILE NOT ENDFILE(MEMORY_FILE) AND I < COUNT - 2 LOOP
            READLINE(MEMORY_FILE, TEXT_LINE);
            I := I + 1;
        END LOOP;

        WHILE NOT ENDFILE(MEMORY_FILE) LOOP
            READLINE(MEMORY_FILE, TEXT_LINE);
            READ(TEXT_LINE, BINARY_TEXT_LINE);
            -- REPORT "TEXT_LINE INSIDE MEMORY LOOP: "& INTEGER'IMAGE(TO_INTEGER(UNSIGNED(TO_STDLOGICVECTOR(BINARY_TEXT_LINE))));
            MEMORY_CONTENT(COUNT) := TO_STDLOGICVECTOR(BINARY_TEXT_LINE);
            COUNT := COUNT + 1;
        END lOOP;

        FILE_CLOSE(MEMORY_FILE);
        RETURN MEMORY_CONTENT;

    END FUNCTION FILL_MEMORY;
    
    SIGNAL INSTRUCTION_MEMORY : MEMORY_TYPE := FILL_MEMORY;

BEGIN
    PROCESS(CLK) IS
        BEGIN
        IF FALLING_EDGE(CLK) THEN
            IF WR = '1' THEN  
                INSTRUCTION_MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))) <= DATA_IN;
            END IF;
            DATA_OUT <= INSTRUCTION_MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)));
        END IF;
    END PROCESS;
END BEHAVIORAL;