library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity controlUnit is port (
Instruction:in std_logic_vector(6 downto 0);
 ALU_SELECTORS:out std_logic_vector(3 downto 0);
 TWO_FETCHES,OP_GROUP:out std_logic_vector(1 downto 0);
 BRANCH,MR,MW,P_IN,P_OUT,SP_INC,SP_DEC,WB1,WB2,CALL,RET,
ALU_ENABLE,RTI,NO_OPERANDS,IGNORE_RSRC2:out std_logic) ;
end controlUnit ;

architecture Behavioral of controlUnit is
begin
process(Instruction)
begin
case (Instruction) is
when "0000000" => --nop
BRANCH <='0';
MR <='0';
MW <='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="00";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='1';
IGNORE_RSRC2 <='1';
when
"0000001" => --not
BRANCH<='0';
ALU_SELECTORS<="0000";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="00";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when
 "0000010" => --inc
BRANCH<='0';
ALU_SELECTORS<="0001";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="00";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "0000011" => --dec
BRANCH<='0';
ALU_SELECTORS<="0010";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="00";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "0000100" => --out
BRANCH<='0';
MR<='0';
MW<='1';
P_IN<='0';
P_OUT<='1';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="00";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';

when
"0000101" => --in
BRANCH<='0';
MR<='1';
MW<='0';
P_IN<='1';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="00";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "0100000" => --jz
BRANCH<='1';
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="01";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "0100001" => --jmp
BRANCH<='0';
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="01";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "0100010" => --call
BRANCH<='0';
MR<='0';
MW<='1';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='1';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="01";
CALL<='1';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "0100111" => --ret
BRANCH<='0';
MR<='1';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='1';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="01";
CALL<='0';
RET<='1';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='1';
IGNORE_RSRC2 <='1';
when "0100101" => --rti
BRANCH<='0';
MR<='1';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='1';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="01";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='1';
NO_OPERANDS <='1';
IGNORE_RSRC2 <='1';
when "1000000" => --swap
BRANCH<='0';
ALU_SELECTORS<="0011";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='1';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='0';
when "1000001" => --add
BRANCH<='0';
ALU_SELECTORS<="0100";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='0';
when "1000010" => --or
 BRANCH<='0';
ALU_SELECTORS<="1000";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='0';
when "1000011" => --sub
 BRANCH<='0';
ALU_SELECTORS<="0110";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='0';
when "1000100" => --and
BRANCH<='0';
ALU_SELECTORS<="0111";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='1';
WB2<='0';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='0';
when "1001101" => --iadd
 BRANCH<='0';
ALU_SELECTORS<="0101";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="01";
WB1<='1';
WB2<='0';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "1001110" => --shl
BRANCH<='0';
ALU_SELECTORS<="1001";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="01";
WB1<='0';
WB2<='1';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "1001111" => --shr
BRANCH<='0';
ALU_SELECTORS<="1011";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="01";
WB1<='0';
WB2<='1';
OP_GROUP<="10";
CALL<='0';
RET<='0';
ALU_ENABLE<='1';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "1100000" => --push
BRANCH<='0';
MR<='0';
MW<='1';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='1';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="11";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "1100001" => --pop
 BRANCH<='0';
MR<='1';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='1';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="11";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "1101010" => --ldm
BRANCH<='0';
MR<='1';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="01";
WB1<='1';
WB2<='0';
OP_GROUP<="11";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "1110101" => --ldd
 BRANCH<='0';
MR<='1';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="10";
WB1<='1';
WB2<='0';
OP_GROUP<="11";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when "1110110" => --std
BRANCH<='0';
MR<='0';
MW<='1';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="10";
WB1<='0';
WB2<='0';
OP_GROUP<="11";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='1';
when others =>
BRANCH<='0';
ALU_SELECTORS<="0000";
MR<='0';
MW<='0';
P_IN<='0';
P_OUT<='0';
SP_INC<='0';
SP_DEC<='0';
TWO_FETCHES<="00";
WB1<='0';
WB2<='0';
OP_GROUP<="00";
CALL<='0';
RET<='0';
ALU_ENABLE<='0';
RTI<='0';
NO_OPERANDS <='0';
IGNORE_RSRC2 <='0';
end case;
end process ;
end Behavioral;
