LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MEMORY_STAGE IS
    PORT (
        -------------------------------- INPUT --------------------------------
        CLK, RST : IN STD_LOGIC;
        EX_MEM_IN : IN STD_LOGIC_VECTOR(111 DOWNTO 0);
        INT : IN STD_LOGIC;
        INSTRUCTION_MEMORY_WR : IN STD_LOGIC;
        CURRENT_PC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        IN_PORT : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        FLAG_REG_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        INSTRUCTION_MEMORY_INPUT : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        INSTRUCTION_MEMORY_ADDRESS : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        -------------------------------- OUTPUT -------------------------------
        DATA_MEMORY_OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        INSTRUCTION_MEMORY_OUTPUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        OUT_PORT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        INTERRUPT_1 : OUT STD_LOGIC;
        RETURN_INT : OUT STD_LOGIC;
        MEM_WB_OUT : OUT STD_LOGIC_VECTOR(72 DOWNTO 0);
        BufferWriteEnable: IN STD_LOGIC 
    );
END MEMORY_STAGE;

ARCHITECTURE DATAFLOW OF MEMORY_STAGE IS
    SIGNAL SP_INCREMENT : STD_LOGIC;
    SIGNAL SP_DECREMENT : STD_LOGIC;
    SIGNAL INTERRUPT_1_SIGNAL : STD_LOGIC;
    SIGNAL INTERRUPT_2 : STD_LOGIC;
    SIGNAL RETURN_INTERRUPT : STD_LOGIC;
    SIGNAL MEMORY_WRITE : STD_LOGIC;
    SIGNAL MEMORY_READ : STD_LOGIC;
    ----------------------- EX/MEM BUFFER INPUT SIGNALS -----------------------
    SIGNAL SP_INC : STD_LOGIC;
    SIGNAL SP_DEC : STD_LOGIC;
    SIGNAL MW : STD_LOGIC;
    SIGNAL MR : STD_LOGIC;
    SIGNAL RTI : STD_LOGIC;
    SIGNAL CALL : STD_LOGIC;
    SIGNAL P_IN : STD_LOGIC;
    SIGNAL P_OUT : STD_LOGIC;
    SIGNAL BUFFER_PC : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL OPERAND_1 : STD_LOGIC_VECTOR (31 DOWNTO 0); -- RESULT
    SIGNAL OPERAND_2 : STD_LOGIC_VECTOR (31 DOWNTO 0); -- EFFECTIVE ADDRESS
    SIGNAL WRITE_REG_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
    SIGNAL WRITE_REG_2 : STD_LOGIC_VECTOR (2 DOWNTO 0);
    ------------------------- MUX TEMP OUTPUT SIGNALS -------------------------
    SIGNAL TEMP_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL TEMP_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL TEMP_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL TEMP_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL TEMP_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL TEMP_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL STACK_POINTER_TEMP : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL CONDITION_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
    SIGNAL CONDITION_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
    ------------------------------ COMPONENTS I/O -----------------------------
    SIGNAL STACK_POINTER_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL STACK_POINTER_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL DATA_MEMORY_DATA_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL DATA_MEMORY_DATA_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL DATA_MEMORY_ADDRESS : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL INSTRUCTION_MEMORY_DATA_OUT : STD_LOGIC_VECTOR (15 DOWNTO 0);
    SIGNAL COMPUTED_OPERAND_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
    SIGNAL MEM_WB_IN : STD_LOGIC_VECTOR (72 DOWNTO 0);


    COMPONENT MEM_WB_BUFFER IS
        PORT (
            CLK, RST, WRITE_ENABLE : IN STD_LOGIC;
            REG_IN : IN STD_LOGIC_VECTOR (72 DOWNTO 0);
            REG_OUT : OUT STD_LOGIC_VECTOR (72 DOWNTO 0));
    END COMPONENT;

    -- STACK REGISTER
    COMPONENT REG IS
        GENERIC (N : INTEGER := 32);
        PORT (
            D : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
            RST, CLK, WR_ENABLE : IN STD_LOGIC;
            Q : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0));
    END COMPONENT;

    COMPONENT DFF IS
        GENERIC (N : INTEGER := 32);
        PORT (
            D : IN STD_LOGIC;
            RST, CLK : IN STD_LOGIC;
            Q : OUT STD_LOGIC
        );
    END COMPONENT;

    COMPONENT INSTRUCTION_MEMORY IS
        GENERIC (
            WORD_SIZE : INTEGER := 16;
            ADDRESS_WIDTH : INTEGER := 32;
            MEMORY_SIZE : INTEGER := 4096);
        PORT (
            WR : IN STD_LOGIC;
            CLK : IN STD_LOGIC;
            ADDRESS : IN STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
            DATA_IN : IN STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
            DATA_OUT : OUT STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0)
        );
    END COMPONENT;

    COMPONENT DATA_MEMORY IS
        GENERIC (
            WORD_SIZE : INTEGER := 16;
            ADDRESS_WIDTH : INTEGER := 32;
            MEMORY_SIZE : INTEGER := 4096);
        PORT (
            WR : IN STD_LOGIC;
            CLK : IN STD_LOGIC;
            ADDRESS : IN STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
            DATA_IN : IN STD_LOGIC_VECTOR(WORD_SIZE * 2 - 1 DOWNTO 0);
            DATA_OUT : OUT STD_LOGIC_VECTOR(WORD_SIZE * 2 - 1 DOWNTO 0)
        );
    END COMPONENT;

BEGIN
    
    MR <= EX_MEM_IN(111);
    MW <= EX_MEM_IN(110);
    P_IN <= EX_MEM_IN(109);
    P_OUT <= EX_MEM_IN(108);
    SP_INC <= EX_MEM_IN(107);
    SP_DEC <= EX_MEM_IN(106);
    CALL <= EX_MEM_IN(103);
    RTI <= EX_MEM_IN(102);
    OPERAND_1 <= EX_MEM_IN(101 DOWNTO 70); -- ALU RESULT
    OPERAND_2 <= EX_MEM_IN(69 DOWNTO 38); -- EFFECTIVE ADDRESS
    BUFFER_PC <= EX_MEM_IN(37 DOWNTO 6);
    WRITE_REG_1 <= EX_MEM_IN(5 DOWNTO 3);
    WRITE_REG_2 <= EX_MEM_IN(2 DOWNTO 0);

    SP_DECREMENT <= INTERRUPT_2 OR INT OR SP_DEC;
    SP_INCREMENT <= RETURN_INTERRUPT OR SP_INC;
    MEMORY_WRITE <= INT OR MW OR INTERRUPT_2;
    MEMORY_READ <= RETURN_INTERRUPT OR MR OR INTERRUPT_1_SIGNAL;

    CONDITION_1 <= SP_INC & SP_DECREMENT;
    CONDITION_2 <= INTERRUPT_1_SIGNAL & RST;

    WITH P_OUT SELECT OUT_PORT <=
        OPERAND_1 WHEN '1',
        (OTHERS => 'Z') WHEN OTHERS;

    WITH CALL SELECT TEMP_1 <=
        BUFFER_PC WHEN '1',
        OPERAND_1 WHEN OTHERS;

    WITH INT SELECT TEMP_2 <=
        CURRENT_PC WHEN '1',
        TEMP_1 WHEN OTHERS;

    WITH INTERRUPT_2 SELECT DATA_MEMORY_DATA_IN <=
        X"0000000" & FLAG_REG_IN WHEN '1',
        TEMP_2 WHEN OTHERS;

    WITH CONDITION_1 SELECT STACK_POINTER_TEMP <=
        STACK_POINTER_OUT WHEN "11",
        STD_LOGIC_VECTOR(UNSIGNED(STACK_POINTER_OUT)) + 2 WHEN "10",
        STD_LOGIC_VECTOR(UNSIGNED(STACK_POINTER_OUT)) - 2 WHEN "01",
        STACK_POINTER_OUT WHEN OTHERS;

    WITH RST SELECT STACK_POINTER_IN <=
        X"000007FF" WHEN '1',
        STACK_POINTER_TEMP WHEN OTHERS;

    WITH SP_INCREMENT SELECT TEMP_3 <=
        STD_LOGIC_VECTOR(UNSIGNED(STACK_POINTER_OUT)) + 2 WHEN '1',
        OPERAND_2 WHEN OTHERS;

    WITH SP_DECREMENT SELECT TEMP_4 <=
        STACK_POINTER_OUT WHEN '1',
        OPERAND_2 WHEN OTHERS;

    WITH MEMORY_READ SELECT TEMP_5 <=
        TEMP_3 WHEN '1',
        TEMP_4 WHEN OTHERS;

    WITH CONDITION_2 SELECT DATA_MEMORY_ADDRESS <=
        X"00000002" WHEN "11",
        X"00000002" WHEN "10",
        X"00000000" WHEN "01",
        TEMP_5 WHEN OTHERS;
    
    WITH MR SELECT TEMP_6 <=
        DATA_MEMORY_DATA_OUT WHEN '1',
        OPERAND_1 WHEN OTHERS;

    WITH P_IN SELECT COMPUTED_OPERAND_1 <=
        IN_PORT WHEN '1',
        TEMP_6 WHEN OTHERS;
    
    ------------------------------ MEM/WB BUFFER ------------------------------

    MEM_WB_IN(0) <= EX_MEM_IN(105); -- WB1
    MEM_WB_IN(1) <= EX_MEM_IN(104); -- WB2
    MEM_WB_IN(2) <= EX_MEM_IN(102); -- RTI
    MEM_WB_IN(34 DOWNTO 3) <= COMPUTED_OPERAND_1; -- OPERAND 1
    MEM_WB_IN(66 DOWNTO 35) <= EX_MEM_IN(69 DOWNTO 38); -- OPERAND 2
    MEM_WB_IN(69 DOWNTO 67) <= EX_MEM_IN(5 DOWNTO 3); -- WRITE_REG_1
    MEM_WB_IN(72 DOWNTO 70) <= EX_MEM_IN(2 DOWNTO 0); -- WRITE_REG_2

    ---------------------------------- OUTPUT ---------------------------------

    DATA_MEMORY_OUTPUT <= DATA_MEMORY_DATA_OUT;
    INSTRUCTION_MEMORY_OUTPUT <= INSTRUCTION_MEMORY_DATA_OUT;
    INTERRUPT_1 <= INTERRUPT_1_SIGNAL;
    RETURN_INT <= RETURN_INTERRUPT;
    
    ------------------------------- PORT MAPPING ------------------------------

    U1 : REG GENERIC MAP(32) PORT MAP(STACK_POINTER_IN, '0', CLK, '1', STACK_POINTER_OUT);
    U2 : DFF PORT MAP(INT, RST, CLK, INTERRUPT_1_SIGNAL);
    U3 : DFF PORT MAP(INTERRUPT_1_SIGNAL, RST, CLK, INTERRUPT_2);
    U4 : DFF PORT MAP(RTI, RST, CLK, RETURN_INTERRUPT);
    U5 : DATA_MEMORY GENERIC MAP(WORD_SIZE => 16, ADDRESS_WIDTH => 32, MEMORY_SIZE => 4096) PORT MAP(MEMORY_WRITE, CLK, DATA_MEMORY_ADDRESS, DATA_MEMORY_DATA_IN, DATA_MEMORY_DATA_OUT);
    U6 : INSTRUCTION_MEMORY GENERIC MAP(WORD_SIZE => 16, ADDRESS_WIDTH => 32, MEMORY_SIZE => 4096) PORT MAP(INSTRUCTION_MEMORY_WR, CLK, INSTRUCTION_MEMORY_ADDRESS, INSTRUCTION_MEMORY_INPUT, INSTRUCTION_MEMORY_DATA_OUT);
    U7 : MEM_WB_BUFFER PORT MAP(CLK, RST, BufferWriteEnable, MEM_WB_IN, MEM_WB_OUT);

END DATAFLOW;