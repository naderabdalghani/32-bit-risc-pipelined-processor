LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY EXECUTIONSTAGE IS
    PORT (
    ID_EX     : IN  STD_LOGIC_VECTOR(129 DOWNTO 0); 
    EX_MEM_IN     : IN  STD_LOGIC_VECTOR(31 DOWNTO 0); 
    MEM_WB     : IN  STD_LOGIC_VECTOR(31 DOWNTO 0); 
    RESET,CLOCK : IN STD_LOGIC ;
    SELFORWARDINGUNIT1  : IN  STD_LOGIC_VECTOR(1 DOWNTO 0); 
    SELFORWARDINGUNIT2  : IN  STD_LOGIC_VECTOR(1 DOWNTO 0); 
    RTIFROMWB : IN STD_LOGIC ;
    CCRFROMWB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    CCR_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    WRONGDECISION : OUT STD_LOGIC ;
    FROM_EXECUTION_STAGE : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    EX_MEM_OUT     : OUT  STD_LOGIC_VECTOR(112 DOWNTO 0);
    BufferWriteEnable : IN STD_LOGIC 
    );
END EXECUTIONSTAGE;

ARCHITECTURE DATAFLOW OF EXECUTIONSTAGE IS
 SIGNAL CHECK1 : STD_LOGIC;
 SIGNAL CHECK2 : STD_LOGIC;
 SIGNAL CHECK3 : STD_LOGIC;
 SIGNAL CHECK4 : STD_LOGIC;
 SIGNAL CCR_ENABLE : STD_LOGIC;
 SIGNAL ALUENABLE : STD_LOGIC;
 SIGNAL SELALU   :  STD_LOGIC_VECTOR(3 DOWNTO 0);
 SIGNAL RESULT1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
 SIGNAL RESULT2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
 SIGNAL OPERAND_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
 SIGNAL OPERAND_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
 SIGNAL CCR_ALU : STD_LOGIC_VECTOR (3 DOWNTO 0);
 SIGNAL CCR_REG : STD_LOGIC_VECTOR (3 DOWNTO 0);
 SIGNAL CCR_REG_INPUT : STD_LOGIC_VECTOR (3 DOWNTO 0);
 SIGNAL BUFF_IN : STD_LOGIC_VECTOR (112 DOWNTO 0);

COMPONENT EX_MEM_BUFFER IS
PORT ( CLOCK, RESET,WRITEENABLE : IN STD_LOGIC;
 REG_IN : IN STD_LOGIC_VECTOR (112 DOWNTO 0);
 REG_OUT : OUT STD_LOGIC_VECTOR (112 DOWNTO 0) );
END COMPONENT; 
COMPONENT ALU IS
  GENERIC ( 
     N: INTEGER := 32  
    );
  
    PORT (
    A, B     : IN  STD_LOGIC_VECTOR(N-1 DOWNTO 0); 
    ENABLE,RESET : IN STD_LOGIC ;
    SEL  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0); 
    RES   : OUT  STD_LOGIC_VECTOR(N-1 DOWNTO 0);
    CCR : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
    );
END COMPONENT; 

COMPONENT CONDITIONCODEREGISTER IS
 PORT ( CLOCK, RESET,WRITEENABLE : IN STD_LOGIC;
 CCRIN : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
 CCROUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0) );
END COMPONENT; 


 BEGIN
 CCR_ENABLE<= ALUENABLE OR RTIFROMWB;
ALUENABLE<= ID_EX(112);
SELALU<= ID_EX(110 DOWNTO 107);
WITH SELFORWARDINGUNIT1 SELECT OPERAND_1 <= -- MUX 1 --
	MEM_WB WHEN "10",
	EX_MEM_IN WHEN "01",
	ID_EX(101 DOWNTO 70) WHEN "00",
	ID_EX(101 DOWNTO 70) WHEN OTHERS;


WITH SELFORWARDINGUNIT2 SELECT OPERAND_2 <= -- MUX 2 --
	MEM_WB WHEN "10",
	EX_MEM_IN WHEN "01",
	ID_EX(69 DOWNTO 38) WHEN "00",
	ID_EX(69 DOWNTO 38) WHEN OTHERS;

WITH SELALU SELECT RESULT2 <= -- MUX 3 -- HANDLING SWAP BY PASSING B IN ALU AND OPERAND ONE GET INTO PLACE OF OPERAND 2 IN BUFFER
        RESULT1 WHEN "1001" | "1011",
        OPERAND_2 WHEN OTHERS;



CHECK1<= ( ID_EX (102) XOR CCR_REG(0) ) AND ID_EX (123) ;
CHECK2<= (NOT(ID_EX (102)) AND NOT(ID_EX (123))) AND CHECK4;
CHECK4<= (NOT (ID_EX (104)) AND ID_EX (103)) AND (NOT (ID_EX (113) OR ID_EX (111)));
CHECK3<= CHECK1 OR CHECK2;
WITH CHECK3 SELECT WRONGDECISION <=
	'1' WHEN '1',
        '0' WHEN OTHERS;

WITH ID_EX (102) SELECT FROM_EXECUTION_STAGE <=
	OPERAND_1 WHEN '0',
	ID_EX(37 DOWNTO 6) WHEN OTHERS;


--HANDLING RTI FROM WB
WITH RTIFROMWB SELECT CCR_REG_INPUT <=
	CCRFROMWB WHEN '1',
        CCR_ALU WHEN OTHERS;

-- OUT 
BUFF_IN (2 DOWNTO 0) <= ID_EX(2 DOWNTO 0);
BUFF_IN (5 DOWNTO 3) <= ID_EX(5 DOWNTO 3);
BUFF_IN (37 DOWNTO 6) <= ID_EX(37 DOWNTO 6);
BUFF_IN (69 DOWNTO 38) <= RESULT2;
BUFF_IN (101 DOWNTO 70) <= RESULT1;
BUFF_IN (102) <= ID_EX(111);
BUFF_IN (111 DOWNTO 103) <= ID_EX(122 DOWNTO 114);
BUFF_IN(112)<= ID_EX(113);
CCR_OUT<=CCR_REG;
-- PORT MAPPING
U1: ALU GENERIC MAP(32)
            PORT MAP(OPERAND_1, OPERAND_2, ID_EX(112),RESET, ID_EX(110 DOWNTO 107),RESULT1,CCR_ALU);
U2: CONDITIONCODEREGISTER  PORT MAP(CLOCK, RESET,CCR_ENABLE ,CCR_REG_INPUT,CCR_REG);
U3: EX_MEM_BUFFER  PORT MAP(CLOCK, RESET,BufferWriteEnable, BUFF_IN,EX_MEM_OUT);

END DATAFLOW;